--
-- VHDL Architecture ece411.Cache_Check.untitled
--
-- Created:
--          by - ravi7.ews (linux-a2.ews.illinois.edu)
--          at - 15:17:47 02/17/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Cache_Check IS
   PORT( 
      clk : IN     std_logic
   );

-- Declarations

END Cache_Check ;

--
ARCHITECTURE untitled OF Cache_Check IS
BEGIN
END ARCHITECTURE untitled;


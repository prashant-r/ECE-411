--
-- VHDL Architecture ece411.SignExt5.untitled
--
-- Created:
--          by - ravi7.ews (gelib-057-36.ews.illinois.edu)
--          at - 15:32:20 01/29/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY SignExt5 IS
   PORT( 
      clk  : IN     std_logic;
      sig0 : IN     std_logic
   );

-- Declarations

END SignExt5 ;

--
ARCHITECTURE untitled OF SignExt5 IS
BEGIN
END ARCHITECTURE untitled;


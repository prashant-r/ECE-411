--
-- VHDL Architecture ece411.ADJ11out.untitled
--
-- Created:
--          by - aikara2.ews (gelib-057-23.ews.illinois.edu)
--          at - 22:53:09 03/17/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY ADJ11out IS
   PORT( 
      RESET_L  : IN     STD_LOGIC;
      clk      : IN     std_logic;
      offset11 : IN     LC3B_offset11;
      adj11out : OUT    LC3b_word
   );

-- Declarations

END ADJ11out ;

--
ARCHITECTURE untitled OF ADJ11out IS
BEGIN
  ADJ11out <= offset11(10) & offset11(10) & offset11(10) & offset11(10) & offset11 & '0' AFTER DELAY_MUX2;
END ARCHITECTURE untitled;



--
-- VHDL Architecture ece411.ByteMux.untitled
--
-- Created:
--          by - ravi7.ews (linux-a1.ews.illinois.edu)
--          at - 14:47:07 02/23/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY ByteMux IS
   PORT( 
      F      : IN     STD_LOGIC;
      High_A : IN     LC3b_BYTE;
      High_b : IN     LC3B_BYTE;
      HighAB : OUT    LC3B_BYTE
   );

-- Declarations

END ByteMux ;

--
ARCHITECTURE untitled OF ByteMux IS
  BEGIN
 PROCESS (High_B, High_A, F)
  variable state : LC3b_byte;
 BEGIN
  case F is
   when '0' =>
  		state := High_a;
			when '1' =>
				state := hIGH_B;
			when others =>
				state := (OTHERS => 'X');
		end case;
		hIGHab <= state after delay_MUX2;
	END PROCESS;
END ARCHITECTURE untitled;


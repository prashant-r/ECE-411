--
-- VHDL Architecture ece411.Word2Byte.untitled
--
-- Created:
--          by - ravi7.ews (linux-a1.ews.illinois.edu)
--          at - 14:53:22 02/23/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Word2Byte IS
   PORT( 
      Potential_word : IN     LC3b_word;
      High_b         : OUT    LC3B_BYTE;
      Low_B          : OUT    LC3B_BYTE
   );

-- Declarations

END Word2Byte ;

--
ARCHITECTURE untitled OF Word2Byte IS
BEGIN
  High_b <= Potential_word( 15 DOWNTO 8);
  Low_b <= Potential_word( 7 DOWNTO 0);
END ARCHITECTURE untitled;


--
-- VHDL Architecture ece411.ZeroGen.untitled
--
-- Created:
--          by - aikara2.ews (gelib-057-38.ews.illinois.edu)
--          at - 20:20:18 03/18/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY ZeroGen IS
   PORT( 
      RESET_L  : IN     STD_LOGIC;
      clk      : IN     std_logic;
      Zero_Out : OUT    LC3b_word
   );

-- Declarations

END ZeroGen ;

--
ARCHITECTURE untitled OF ZeroGen IS
BEGIN
  
  Zero_Out <= "0000000000000000" after delay_reg; 
  
END ARCHITECTURE untitled;


--
-- VHDL Architecture ece411.Sure00.untitled
--
-- Created:
--          by - ravi7.ews (linux-a1.ews.illinois.edu)
--          at - 12:50:58 03/23/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Sure00 IS
   PORT( 
      clk      : IN     std_logic;
      zerozero : OUT    std_logic_vector (1 DOWNTO 0)
   );

-- Declarations

END Sure00 ;

--
ARCHITECTURE untitled OF Sure00 IS
BEGIN
  zerozero <= "00";
END ARCHITECTURE untitled;

